module dmemory #()
(
    
);



endmodule
